`ifndef _PC_REG_V_
`define _PC_REG_V_

// 1. 程序计数器模块接口部分：
module pc_reg( // 时序电路
    input wire      clk, // 声明了一个名为clk的输入端口，类型为wire。这是时钟信号，用于同步电路操作，控制PC寄存器的更新时机。
    input wire      rst, // 声明了一个名为rst的输入端口，类型为wire。这是复位信号，用于重置PC寄存器(通常是0)。
    input wire[31:0] jump_addr_i,
    input wire      jump_en_i,    
    // [31:0] 是Verilog中的位宽描述符，表示一个32位的数据信号或变量。这种表示方法指定了位的范围：
        // 31是最高位(Most Significant Bit, MSB)
        // 0是最低位(Least Significant Bit, LSB)
        // 总共有32位(从0到31，包含0和31)
    output reg[31:0] pc_o // 声明了一个名为pc_o的输出端口，是32位宽的寄存器类型变量，作为输出端口，用来存储当前指令地址。
);  

// 补充：
// wire 类型：在Verilog中，wire 是一种数据类型，表示电路中的物理连线。它的特点是：
    // 不存储值，只传递值
    // 连接模块之间或模块内部不同部件的信号
    // 不能在过程块中(如always块)被赋值
    // 代表组合逻辑中的连接
// 简单来说，wire 就像电路图中的导线，它可以传递信号，但不能存储信号。



// 2. 功能实现部分：
    // 这定义了一个时序逻辑块，只在时钟信号(clk)的上升沿触发。意味着以下代码块中的操作只会在时钟从0变为1的瞬间执行。
    always @(posedge clk) begin 
             
        // 1) 查复位信号(rst)是否为低电平(0)。
        // 2) rst == 1'b0使用二进制('b)是因为：
            // 复位信号通常是一个单一位的控制信号
            // 1'b0明确表示一个1位的二进制0
            // 对于单位的控制信号和标志位，通常习惯使用二进制表示
        if(rst == 1'b0) 
            // 如果复位信号有效(为0)，则将PC寄存器地址值重置为0。32'b0表示32位的二进制0，<=是非阻塞赋值运算符，
            // 在 always @(posedge clk) 块内，适用于时序逻辑。
            pc_o <= 32'b0;
        else if(jump_en_i == 1'b1)
            pc_o <= jump_addr_i;
        else
            // 如果复位信号无效(为1)，则PC寄存器的值增加4。32'd4表示32位的十进制值4。PC增加4是因为在大多数32位架构中，每条指令占4个字节(32位)。
            pc_o <= pc_o + 32'd4;
    end

// 补充：
// 时序逻辑（如 always @posedge clk 块）中应该使用非阻塞赋值 <=，原因是：
    // 它模拟了硬件中寄存器的实际行为（同时更新）
    // 避免了由于赋值顺序导致的竞争条件
    // 确保模拟结果与实际硬件行为一致
// 1. 使用<=（非阻塞赋值）时机：
    // 1) 在时序逻辑中：所有由时钟控制的always块中
    // 2) 描述寄存器行为时：任何需要存储状态的电路元件
    // 3) 同步电路设计中：所有触发器和寄存器更新
// 2. 使用=（阻塞赋值）时机：
    // 1) 在组合逻辑中：对应于纯组合电路的always块
    // 2) 临时变量赋值：在过程块中使用的中间变量
    // 3) 初始化块中
// 总结：时钟相关使用 <=，组合逻辑使用 =。

endmodule
`endif