`ifndef _ROM_V_
`define _ROM_V_
module rom(
    input wire[31:0] inst_addr_i,
    output reg[31:0] inst_o
);

// 补充：reg vs. wire
// 什么时候用 reg？
    // 当信号在 always 块中被赋值（即过程性赋值）。
    // 作为 output 时，如果它是 always 块内的变量。
// 什么时候用 wire？
    // 当信号用 assign 赋值（连续赋值）。
    // 作为 input 时（因为 input 默认是 wire）。
    // 作为 output 时，如果它直接连接到 assign 或者是子模块的 wire。
// 简易判断法则：
    // 如果信号在always块中被赋值 → 使用reg
    // 如果信号通过assign语句赋值 → 使用wire
    // 所有模块输入必须是wire   
    // 模块输出可以是reg或wire，取决于它如何被赋值



    reg[31:0] rom_mem[0:4095]; // 4096 个 32'b的空间

    // 内存地址与指令的关系：
        // 字节地址:   0   1   2   3   4   5   6   7   8   9  10  11
        //            |---|---|---|---|---|---|---|---|---|---|---|---|
        // 指令编号:   |    指令0     |    指令1     |    指令2     |
        // 现在，如果我要访问指令1，我需要提供地址4。但ROM数组的索引不是按字节地址存储的，而是按指令编号：
        // Copyrom_mem[0] = 指令0的内容
        // rom_mem[1] = 指令1的内容
        // rom_mem[2] = 指令2的内容
        // 因此需要将字节地址转换为指令编号。转换公式是：
        // Copy指令编号 = 字节地址 ÷ 4
        // 在二进制中，除以4等同于右移2位。例如：

        // 10进制的8，二进制是1000
        // 右移2位后变成10 (二进制)，等于10进制的2
        // 8 ÷ 4 = 2
        // 所以，inst_addr_i>>2就是把指令的字节地址转换为ROM数组中的索引位置。
        // 例如：
        // 当CPU请求一条32位指令时，它提供的是这条指令的起始字节地址。
        // 如果CPU请求地址4，4>>2 = 1，就会返回rom_mem[1]的内容
        // 如果CPU请求地址8，8>>2 = 2，就会返回rom_mem[2]的内容
        // 这就是为什么需要右移2位(>>2)，它把字节地址转换为指令的索引位置。
            // 二进制右移（>>）是将所有位向右移动指定的位数，最左边添加0（对于无符号数）。这相当于除以2的n次方，其中n是右移的位数。
                // 例如，对于二进制数 1010（十进制10）：
                // 右移1位：1010 >> 1 = 0101（十进制5）
                // 右移2位：1010 >> 2 = 0010（十进制2）
                // 右移3位：1010 >> 3 = 0001（十进制1）
            // 左移操作（<<）正好与右移相反，它将所有二进制位向左移动指定的位数，右边补0。左移相当于乘以2的n次方，其中n是左移的位数。
    always @(*)begin
            inst_o = rom_mem[inst_addr_i>>2];
        end

endmodule
`endif